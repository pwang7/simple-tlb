`include "sample_tests.vh"
else if(testname =="bypass_test")
begin
    // Since the main logic is in mkXDMATestbench, there is left empty.
end
